
module top_module(
    output one
);

    // Always assign the output to 1 (logic high)
    assign one = 1'b1;

endmodule
