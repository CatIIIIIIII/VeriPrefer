
module top_module(
    input in,
    output out
);
    // Assign the output port to the same value as the input port
    assign out = in;
endmodule
