
module top_module(
    output zero
);

    // Assign the output zero to a constant value of 0
    assign zero = 1'b0;

endmodule
