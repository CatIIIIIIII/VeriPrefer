
module top_module(
    output zero
);

    // Always assign the output to 0
    assign zero = 0;

endmodule
