
module top_module (
    input [1023:0] in,
    input [7:0] sel,
    output [3:0] out
);

always @(*) begin
    case (sel)
        8'b00000000: out = in[3:0];
        8'b00000001: out = in[7:4];
        8'b00000010: out = in[11:8];
        8'b00000011: out = in[15:12];
        8'b00000100: out = in[19:16];
        8'b00000101: out = in[23:20];
        8'b00000110: out = in[27:24];
        8'b00000111: out = in[31:28];
        8'b00001000: out = in[35:32];
        8'b00001001: out = in[39:36];
        8'b00001010: out = in[43:40];
        8'b00001011: out = in[47:44];
        8'b00001100: out = in[51:48];
        8'b00001101: out = in[55:52];
        8'b00001110: out = in[59:56];
        8'b00001111: out = in[63:60];
        8'b00010000: out = in[67:64];
        8'b00010001: out = in[71:68];
        8'b00010010: out = in[75:72];
        8'b00010011: out = in[79:76];
        8'b00010100: out = in[83:80];
        8'b00010101: out = in[87:84];
        8'b00010110: out = in[91:88];
        8'b00010111: out = in[95:92];
        8'b00011000: out = in[99:96];
        8'b00011001: out = in[103:100];
        8'b00011010: out = in[107:104];
        8'b00011011: out = in[111:108];
        8'b00011100: out = in[115:112];
        8'b00011101: out = in[119:116];
        8'b00011110: out = in[123:120];
        8'b00011111: out = in[127:124];
        8'b00100000: out = in[131:128];
        8'b00100001: out = in[135:132];
        8'b00100010: out = in[139:136];
        8'b00100011: out = in[143:140];
        8'b00100100: out = in[147:144];
        8'b00100101: out = in[151:148];
        8'b00100110: out = in[155:152];
        8'b00100111: out = in[159:156];
        8'b00101000: out = in[163:160];
        8'b00101001: out = in[167:164];
        8'b00101010: out = in[171:168];
        8'b00101011: out = in[175:172];
        8'b00101100: out = in[179:176];
        8'b00101101: out = in[183:180];
        8'b00101110: out = in[187:184];
        8'b00101111: out = in[191:188];
        8'b00110000: out = in[195:192];
        8'b00110001: out = in[199:196];
        8'b00110010: out = in[203:200];
        8'b00110011: out = in[207:204];
        8'b00110100: out = in[211:208];
        8'b00110101: out = in[215:212];
        8'b00110110: out = in[219:216];
        8'b00110111: out = in[223:220];
        8'b00111000: out = in[227:224];
        8'b00111001: out = in[231:228];
        8'b00111010: out = in[235:232];
        8'b00111011: out = in[239:236];
        8'b00111100: out = in[243:240];
        8'b00111101: out = in[247:244];
        8'b00111110: out = in[251:248];
        8'b00111111: out = in[255:252];
        8'b01000000: out = in[259:256];
        8'b01000001: out = in[263:260];
        8'b01000010: out = in[267:264];
        8'b01000011: out = in[271:268];
        8'b01000100: out = in[275:272];
        8'b01000101: out = in[279:276];
        8'b01000110: out = in[283:280];
        8'b01000111: out = in[287:284];
        8'b01001000: out = in[291:288];
        8'b01001001: out = in[295:292];
        8'b01001010: out = in[299:296];
        8'b01001011: out = in[303:300];
        8'b01001100: out = in[307:304];
        8'b01001101: out = in[311:308];
        8'b01001110: out = in[315:312];
        8'b01001111: out = in[319:316];
        8'b01010000: out = in[323:320];
        8'b01010001: out = in[327:324];
        8'b01010010: out = in[331:328];
        8'b01010011: out = in[335:332];
        8'b01010100: out = in[339:336];
        8'b01010101: out = in[343:340];
        8'b01010110: out = in[347:344];
        8'b01010111: out = in[351:348];
        8'b01011000: out = in[355:352];
        8'b01011001: out = in[359:356];
        8'b01011010: out = in[363:360];
        8'b01011011: out = in[367:364];
        8'b01011100: out = in[371:368];
        8'b01011101: out = in[375:372];
        8'b01011110: out = in[379:376];
        8'b01011111: out = in[383:380];
        8'b01100000: out = in[387:384];
        8'b01100001: out = in[391:388];
        8'b01100010: out = in[395:392];
        8'b01100011: out = in[399:396];
        8'b01100100: out = in[403:400];
        8'b01100101: out = in[407:404];
        8'b01100110: out = in[411:408];
        8'b01100111: out = in[415:412];
        8'b01101000: out = in[419:416];
        8'b01101001: out = in[423:420];
        8'b01101010: out = in[427:424];
        8'b01101011: out = in[431:428];
        8'b01101100: out = in[435:432];
        8'b01101101: out = in[439:436];
        8'b01101110: out = in[443:440];
        8'b01101111: out = in[447:444];
        8'b01110000: out = in[451:448];
        8'b01110001: out = in[455:452];
        8'b01110010: out = in[459:456];
        8'b01110011: out = in[463:460];
        8'b01110100: out = in[467:464];
        8'b01110101: out = in[471:468];
        8'b01110110: out = in[475:472];
        8'b01110111: out = in[479:476];
        8'b01111000: out = in[483:480];
        8'b01111001: out = in[487:484];
        8'b01111010: out = in[491:488];
        8'b01111011: out = in[495:492];
        8'b01111100: out = in[499:496];
        8'b01111101: out = in[503:500];
        8'b01111110: out = in[507:504];
        8'b01111111: out = in[511:508];
        8'b10000000: out = in[515:512];
        8'b10000001: out = in[519:516];
        8'b10000010: out = in[523:520];
        8'b10000011: out = in[527:524];
        8'b10000100: out = in[531:528];
        8'b10000101: out = in[535:532];
        8'b10000110: out = in[539:536];
        8'b10000111: out = in[543:540];
        8'b10001000: out = in[547:544];
        8'b10001001: out = in[551:548];
        8'b10001010: out = in[555:552];
        8'b10001011: out = in[559:556];
        8'b10001100: out = in[563:560];
        8'b10001101: out = in[567:564];
        8'b10001110: out = in[571:568];
        8'b10001111: out = in[575:572];
        8'b10010000: out = in[579:576];
        8'b10010001: out = in[583:580];
        8'b10010010: out = in[587:584];
        8'b10010011: out = in[591:588];
        8'b10010100: out = in[595:592];
        8'b10010101: out = in[599:596];
        8'b10010110: out = in[603:600];
        8'b10010111: out = in[607:604];
        8'b10011000: out = in[611:608];
        8'b10011001: out = in[615:612];
        8'b10011010: out = in[619:616];
        8'b10011011: out