`timescale 1 ps/1 ps
`define OK 12
`define INCORRECT 13
module reference_module(
	output one);
	
	assign one = 1'b1;
	
endmodule


module stimulus_gen (
	input clk,
	output reg[511:0] wavedrom_title,
	output reg wavedrom_enable
);


// Add two ports to module stimulus_gen:
//    output [511:0] wavedrom_title
//    output reg wavedrom_enable

	task wavedrom_start(input[511:0] title = "");
	endtask
	
	task wavedrom_stop;
		#1;
	endtask	



	initial begin
		wavedrom_start("Output should be 1");
		repeat(20) @(posedge clk, negedge clk);
		wavedrom_stop();
		
		#1 $finish;
	end
	
endmodule

module testbench;

	typedef struct packed {
		int errors;
		int errortime;
		int errors_one;
		int errortime_one;

		int clocks;
	} stats;
	
	stats stats1;
	
	
	wire[511:0] wavedrom_title;
	wire wavedrom_enable;
	int wavedrom_hide_after_time;
	
	reg clk=0;
	initial forever
		#5 clk = ~clk;

	logic one_ref;
	logic one_dut;

	initial begin 
		$dumpfile("wave.vcd");
		$dumpvars(1, stim1.clk, tb_mismatch ,one_ref,one_dut );
	end


	wire tb_match;		// Verification
	wire tb_mismatch = ~tb_match;
	
	stimulus_gen stim1 (
		.clk,
		.*  );
	reference_module good1 (
		.one(one_ref) );
		
	top_module top_module1 (
		.one(one_dut) );

	
	bit strobe = 0;
	task wait_for_end_of_timestep;
		repeat(5) begin
			strobe <= !strobe;  // Try to delay until the very end of the time step.
			@(strobe);
		end
	endtask	

	
	final begin
		if (stats1.errors_one) $display("Hint: Output '%s' has %0d mismatches. First mismatch occurred at time %0d.", "one", stats1.errors_one, stats1.errortime_one);
		else $display("Hint: Output '%s' has no mismatches.", "one");

		if (stats1.errors == 0) begin
			$display("Your Design Passed");
		end else begin
			$display("Your Design Failed");
		end
		$display("Simulation finished at %0d ps", $time);
		$display("Mismatches: %1d in %1d samples", stats1.errors, stats1.clocks);
	end
	
	// Verification: XORs on the right makes any X in good_vector match anything, but X in dut_vector will only match X.
	assign tb_match = ( { one_ref } === ( { one_ref } ^ { one_dut } ^ { one_ref } ) );
	// Use explicit sensitivity list here. @(*) causes NetProc::nex_input() to be called when trying to compute
	// the sensitivity list of the @(strobe) process, which isn't implemented.
	always @(posedge clk, negedge clk) begin

		stats1.clocks++;
		if (!tb_match) begin
			if (stats1.errors == 0) stats1.errortime = $time;
			stats1.errors++;
		end
		if (one_ref !== ( one_ref ^ one_dut ^ one_ref ))
		begin if (stats1.errors_one == 0) stats1.errortime_one = $time;
			stats1.errors_one = stats1.errors_one+1'b1; end

	end
endmodule
