
module top_module(
    input a, 
    input b,
    output out
);
    // AND gate logic
    assign out = a & b;
endmodule
