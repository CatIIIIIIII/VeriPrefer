
module top_module(
    output out
);

    // Always assign the output to 0
    assign out = 0;

endmodule
