
module top_module(
	input in,
	output out
);

	// NOT gate implementation
	assign out = ~in;

endmodule
