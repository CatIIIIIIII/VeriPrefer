
module top_module(
    input a, 
    input b,
    output out
);
    // Logical AND operation
    assign out = a & b;
endmodule
