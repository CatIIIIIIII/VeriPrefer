
module top_module (
    input a,
    input b,
    input c,
    output w,
    output x,
    output y,
    output z  
);

    // Assigning the values of inputs to outputs
    assign w = a;
    assign x = b;
    assign y = b;
    assign z = c;

endmodule
