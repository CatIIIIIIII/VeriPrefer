
module top_module (
    input [255:0] in,
    input [7:0] sel,
    output out
);

assign out = (sel == 8'd0) ? in[0] :
            (sel == 8'd1) ? in[1] :
            (sel == 8'd2) ? in[2] :
            (sel == 8'd3) ? in[3] :
            (sel == 8'd4) ? in[4] :
            (sel == 8'd5) ? in[5] :
            (sel == 8'd6) ? in[6] :
            (sel == 8'd7) ? in[7] :
            (sel == 8'd8) ? in[8] :
            (sel == 8'd9) ? in[9] :
            (sel == 8'd10) ? in[10] :
            (sel == 8'd11) ? in[11] :
            (sel == 8'd12) ? in[12] :
            (sel == 8'd13) ? in[13] :
            (sel == 8'd14) ? in[14] :
            (sel == 8'd15) ? in[15] :
            (sel == 8'd16) ? in[16] :
            (sel == 8'd17) ? in[17] :
            (sel == 8'd18) ? in[18] :
            (sel == 8'd19) ? in[19] :
            (sel == 8'd20) ? in[20] :
            (sel == 8'd21) ? in[21] :
            (sel == 8'd22) ? in[22] :
            (sel == 8'd23) ? in[23] :
            (sel == 8'd24) ? in[24] :
            (sel == 8'd25) ? in[25] :
            (sel == 8'd26) ? in[26] :
            (sel == 8'd27) ? in[27] :
            (sel == 8'd28) ? in[28] :
            (sel == 8'd29) ? in[29] :
            (sel == 8'd30) ? in[30] :
            (sel == 8'd31) ? in[31] :
            (sel == 8'd32) ? in[32] :
            (sel == 8'd33) ? in[33] :
            (sel == 8'd34) ? in[34] :
            (sel == 8'd35) ? in[35] :
            (sel == 8'd36) ? in[36] :
            (sel == 8'd37) ? in[37] :
            (sel == 8'd38) ? in[38] :
            (sel == 8'd39) ? in[39] :
            (sel == 8'd40) ? in[40] :
            (sel == 8'd41) ? in[41] :
            (sel == 8'd42) ? in[42] :
            (sel == 8'd43) ? in[43] :
            (sel == 8'd44) ? in[44] :
            (sel == 8'd45) ? in[45] :
            (sel == 8'd46) ? in[46] :
            (sel == 8'd47) ? in[47] :
            (sel == 8'd48) ? in[48] :
            (sel == 8'd49) ? in[49] :
            (sel == 8'd50) ? in[50] :
            (sel == 8'd51) ? in[51] :
            (sel == 8'd52) ? in[52] :
            (sel == 8'd53) ? in[53] :
            (sel == 8'd54) ? in[54] :
            (sel == 8'd55) ? in[55] :
            (sel == 8'd56) ? in[56] :
            (sel == 8'd57) ? in[57] :
            (sel == 8'd58) ? in[58] :
            (sel == 8'd59) ? in[59] :
            (sel == 8'd60) ? in[60] :
            (sel == 8'd61) ? in[61] :
            (sel == 8'd62) ? in[62] :
            (sel == 8'd63) ? in[63] :
            (sel == 8'd64) ? in[64] :
            (sel == 8'd65) ? in[65] :
            (sel == 8'd66) ? in[66] :
            (sel == 8'd67) ? in[67] :
            (sel == 8'd68) ? in[68] :
            (sel == 8'd69) ? in[69] :
            (sel == 8'd70) ? in[70] :
            (sel == 8'd71) ? in[71] :
            (sel == 8'd72) ? in[72] :
            (sel == 8'd73) ? in[73] :
            (sel == 8'd74) ? in[74] :
            (sel == 8'd75) ? in[75] :
            (sel == 8'd76) ? in[76] :
            (sel == 8'd77) ? in[77] :
            (sel == 8'd78) ? in[78] :
            (sel == 8'd79) ? in[79] :
            (sel == 8'd80) ? in[80] :
            (sel == 8'd81) ? in[81] :
            (sel == 8'd82) ? in[82] :
            (sel == 8'd83) ? in[83] :
            (sel == 8'd84) ? in[84] :
            (sel == 8'd85) ? in[85] :
            (sel == 8'd86) ? in[86] :
            (sel == 8'd87) ? in[87] :
            (sel == 8'd88) ? in[88] :
            (sel == 8'd89) ? in[89] :
            (sel == 8'd90) ? in[90] :
            (sel == 8'd91) ? in[91] :
            (sel == 8'd92) ? in[92] :
            (sel == 8'd93) ? in[93] :
            (sel == 8'd94) ? in[94] :
            (sel == 8'd95) ? in[95] :
            (sel == 8'd96) ? in[96] :
            (sel == 8'd97) ? in[97] :
            (sel == 8'd98) ? in[98] :
            (sel == 8'd99) ? in[99] :
            (sel == 8'd100) ? in[100] :
            (sel == 8'd101) ? in[101] :
            (sel == 8'd102) ? in[102] :
            (sel == 8'd103) ? in[103] :
            (sel == 8'd104) ? in[104] :
            (sel == 8'd105) ? in[105] :
            (sel == 8'd106) ? in[106] :
            (sel == 8'd107) ? in[107] :
            (sel == 8'd108) ? in[108] :
            (sel == 8'd109) ? in[109] :
            (sel == 8'd110) ? in[110] :
            (sel == 8'd111) ? in[111] :
            (sel == 8'd112) ? in[112] :
            (sel == 8'd113) ? in[113] :
            (sel == 8'd114) ? in[114] :
            (sel == 8'd115) ? in[115] :
            (sel == 8'd116) ? in[116] :
            (sel == 8'd117) ? in[117] :
            (sel == 8'd118) ? in[118] :
            (sel == 8'd119) ? in[119] :
            (sel == 8'd120) ? in[120] :
            (sel == 8'd121) ? in[121] :
            (sel == 8'd122) ? in[122] :
            (sel == 8'd123) ? in[123] :
            (sel == 8'd124) ? in[124] :
            (sel == 8'd125) ? in[125] :
            (sel == 8'd126) ? in[126] :
            (sel == 8'd127) ? in[127] :
            (sel == 8'd128) ? in[128] :
            (sel == 8'd129) ? in[129] :
            (sel == 8'd130) ? in[130] :
            (sel == 8'd131) ? in[131] :
            (sel == 8'd132) ? in[132] :
            (sel == 8'd133) ? in[133] :
            (sel == 8'd134) ? in[134] :
            (sel == 8'd135) ? in[135] :
            (sel == 8'd136) ? in[136] :
            (sel == 8'd137) ? in[137] :
            (sel == 8'd138) ? in[138] :
            (sel == 8'd139) ? in[139] :
            (sel == 8'd140) ? in[140] :
            (sel == 8'd141) ? in[141] :
            (sel == 8'd142) ? in[142] :
            (sel == 8'd143) ? in[143] :
            (sel == 8'd144) ? in[144] :
            (sel == 8'd145) ? in[145] :
            (sel == 8'd146) ? in[146] :
            (sel == 8'd147) ? in[147] :
            (sel == 8'd148) ? in[148] :
            (sel == 8'd149) ? in[149] :
            (sel == 8'd150) ? in[150] :
            (sel == 8'd151) ? in[151] :
            (sel == 8'd152) ? in[152] :
            (sel == 8'd153) ? in[153] :
            (sel == 8'd154) ? in[154] :
            (sel == 8'd155) ? in[155] :
            (sel == 8'd156) ? in[156] :
            (sel == 8'd157) ? in[157] :
            (sel == 8'd158) ? in[158] :
            (sel == 8'd159) ? in[159] :
            (sel == 8'd160) ? in[160] :
            (sel == 8'd161) ? in[161] :
            (sel == 8'd162) ? in[162] :
            (sel == 8'd163) ? in[163] :
            (sel == 8'd164) ? in[164] :
            (sel == 8'd165) ? in[165] :
            (sel == 8'd166) ? in[166] :
            (sel == 8'd167) ? in[167] :
            (sel == 8'd168) ? in[168] :
            (sel == 8'd169) ? in[169] :
            (sel == 8'd170) ? in[170] :
            (sel == 8'd171) ? in[171] :
            (sel == 8'd172) ? in[172] :
            (sel == 8'd173) ? in[173] :
            (sel == 8'd174) ? in[174] :
            (sel == 8'd175) ? in[175] :
            (sel == 8'd176) ? in[176] :
            (sel == 8'd177) ? in[177] :
            (sel == 8'd178) ? in[178] :
            (sel == 8'd179) ? in[179] :
            (sel == 8'd180) ? in[180] :
            (sel == 8'd181) ? in[181] :
            (sel == 8'd182) ? in[182] :
            (sel == 8'd183) ? in[183] :
            (sel == 8'd184) ? in[184] :
            (sel == 8'd185) ? in[185] :
            (sel == 8'd186) ? in[186] :
            (sel == 8'd187) ? in[187] :
            (sel == 8'd188) ? in[188] :
            (sel == 8'd189) ? in[189] :
            (sel == 8'd190) ? in[190] :
            (sel == 8'd191) ? in[191] :
            (sel == 8'd192) ? in[192] :
            (sel == 8'd193) ? in[193] :
            (sel == 8'd194) ? in[194] :
            (sel == 8'd195) ? in[195] :
            (sel == 8'd196) ? in[196] :
            (sel == 8'd197) ? in[197] :
            (sel == 8'd198) ? in[198] :
            (sel == 8'd199) ? in[199] :
            (sel == 8'd200) ? in[200] :
            (sel == 8'd201) ? in[201] :
            (sel == 8'd202) ? in[202] :
            (sel == 8'd203) ? in[203] :
            (sel == 8'd204) ? in[204] :
            (sel == 8'd205) ? in[205] :
            (sel == 8'd206) ? in[206] :
            (sel == 8'd207) ? in[207] :
            (sel == 8'd208) ? in[208] :
            (sel == 8'd209) ? in[209] :
            (sel == 8'd210) ? in[210] :
            (sel == 8'd211) ? in[211] :
            (sel == 8'd212) ? in[212] :
            (sel == 8'd213) ? in[213] :
            (sel == 8'd214) ? in[214] :
            (sel == 8'd