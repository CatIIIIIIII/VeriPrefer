
module top_module (
    input a, 
    input b, 
    output q
);
    // Perform the AND operation between inputs a and b
    assign q = a & b;
endmodule
