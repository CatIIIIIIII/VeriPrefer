
module top_module(
    output one
);

    // Assign the output one to a constant value of 1'b1
    assign one = 1'b1;

endmodule
