
module top_module (
    input a, 
    input b, 
    output q
);
    // Implementing the AND gate
    assign q = a & b;
endmodule
