
module top_module(
    output out
);

    // Assign the output port to a constant value of 0
    assign out = 1'b0;

endmodule
