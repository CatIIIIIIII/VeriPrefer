
module top_module(
    input in,
    output out
);
    // The output is directly assigned the value of the input
    assign out = in;
endmodule
