
module top_module (
    input a,
    input b,
    input c,
    output w,
    output x,
    output y,
    output z
);

// Assigning inputs to outputs as specified
assign w = a;
assign x = b;
assign y = b;
assign z = c;

endmodule
