`timescale 1 ps/1 ps
`define OK 12
`define INCORRECT 13
module reference_module (
	input [2:0] sel,
	input [3:0] data0,
	input [3:0] data1,
	input [3:0] data2,
	input [3:0] data3,
	input [3:0] data4,
	input [3:0] data5,
	output reg [3:0] out
);

	always @(*) begin
		case (sel)
			3'h0: out = data0;
			3'h1: out = data1;
			3'h2: out = data2;
			3'h3: out = data3;
			3'h4: out = data4;
			3'h5: out = data5;
			default: out = 4'b0;
		endcase
	end
	
endmodule


module stimulus_gen (
	input clk,
	output logic [2:0] sel, 
	output logic [3:0] data0,
	output logic [3:0] data1,
	output logic [3:0] data2,
	output logic [3:0] data3,
	output logic [3:0] data4,
	output logic [3:0] data5,
	output reg[511:0] wavedrom_title,
	output reg wavedrom_enable	
);


// Add two ports to module stimulus_gen:
//    output [511:0] wavedrom_title
//    output reg wavedrom_enable

	task wavedrom_start(input[511:0] title = "");
	endtask
	
	task wavedrom_stop;
		#1;
	endtask	



	initial begin
		data0 <= 4'ha;
		data1 <= 4'hb;
		data2 <= 4'hc;
		data3 <= 4'hd;
		data4 <= 4'he;
		data5 <= 4'hf;
		{sel} <= 3'b111;
		@(negedge clk) wavedrom_start("<b>Sel</b> chooses one of the data inputs");
			repeat(8) @(posedge clk) sel <= sel + 1;
		@(negedge clk) wavedrom_stop();

		repeat(100) @(posedge clk, negedge clk) begin
			{data0, data1, data2, data3} <= $urandom;
			{data4, data5, sel} <= $urandom;
		end
		$finish;
	end
	
endmodule

module testbench;

	typedef struct packed {
		int errors;
		int errortime;
		int errors_out;
		int errortime_out;

		int clocks;
	} stats;
	
	stats stats1;
	
	
	wire[511:0] wavedrom_title;
	wire wavedrom_enable;
	int wavedrom_hide_after_time;
	
	reg clk=0;
	initial forever
		#5 clk = ~clk;

	logic [2:0] sel;
	logic [3:0] data0;
	logic [3:0] data1;
	logic [3:0] data2;
	logic [3:0] data3;
	logic [3:0] data4;
	logic [3:0] data5;
	logic [3:0] out_ref;
	logic [3:0] out_dut;

	initial begin 
		$dumpfile("wave.vcd");
		$dumpvars(1, stim1.clk, tb_mismatch ,sel,data0,data1,data2,data3,data4,data5,out_ref,out_dut );
	end


	wire tb_match;		// Verification
	wire tb_mismatch = ~tb_match;
	
	stimulus_gen stim1 (
		.clk,
		.* ,
		.sel,
		.data0,
		.data1,
		.data2,
		.data3,
		.data4,
		.data5 );
	reference_module good1 (
		.sel,
		.data0,
		.data1,
		.data2,
		.data3,
		.data4,
		.data5,
		.out(out_ref) );
		
	top_module top_module1 (
		.sel,
		.data0,
		.data1,
		.data2,
		.data3,
		.data4,
		.data5,
		.out(out_dut) );

	
	bit strobe = 0;
	task wait_for_end_of_timestep;
		repeat(5) begin
			strobe <= !strobe;  // Try to delay until the very end of the time step.
			@(strobe);
		end
	endtask	

	
	final begin
		if (stats1.errors_out) $display("Hint: Output '%s' has %0d mismatches. First mismatch occurred at time %0d.", "out", stats1.errors_out, stats1.errortime_out);
		else $display("Hint: Output '%s' has no mismatches.", "out");

		if (stats1.errors == 0) begin
			$display("Your Design Passed");
		end else begin
			$display("Your Design Failed");
		end
		$display("Simulation finished at %0d ps", $time);
		$display("Mismatches: %1d in %1d samples", stats1.errors, stats1.clocks);
	end
	
	// Verification: XORs on the right makes any X in good_vector match anything, but X in dut_vector will only match X.
	assign tb_match = ( { out_ref } === ( { out_ref } ^ { out_dut } ^ { out_ref } ) );
	// Use explicit sensitivity list here. @(*) causes NetProc::nex_input() to be called when trying to compute
	// the sensitivity list of the @(strobe) process, which isn't implemented.
	always @(posedge clk, negedge clk) begin

		stats1.clocks++;
		if (!tb_match) begin
			if (stats1.errors == 0) stats1.errortime = $time;
			stats1.errors++;
		end
		if (out_ref !== ( out_ref ^ out_dut ^ out_ref ))
		begin if (stats1.errors_out == 0) stats1.errortime_out = $time;
			stats1.errors_out = stats1.errors_out+1'b1; end

	end
endmodule
